module cpu_regfile (
    input logic clk,
    input logic rst_n,
    output logic
);

logic[31:0] registers[31:0];

endmodule