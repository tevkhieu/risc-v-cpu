/*
 ==============================================================================
 Filename  : cpu_top.sv
 Project   : risc-v-cpu
 Author    : Tévchhorpoan Khieu
 Created   : 2025-11-16

 Description:
    - Top-level CPU module definition.

 Notes:
    - WIP
 ==============================================================================
*/

module cpu_top (
    input logic clk,
    input logic rst_n
);
    
endmodule